module Adder(cin,a,b,s,overflow);        
           input[31:0]a;
           input[31:0]b;
           input cin;
           output[31:0]s;
           output overflow;
           wire [30:0]c;
full_adder a1(.Co(c[0]),.S(s[0]),.X(a[0]),.Y(b[0]),.Ci(cin));
full_adder a2(.Co(c[1]),.S(s[1]),.X(a[1]),.Y(b[1]),.Ci(c[0]));
full_adder a3(.Co(c[2]),.S(s[2]),.X(a[2]),.Y(b[2]),.Ci(c[1]));
full_adder a4(.Co(c[3]),.S(s[3]),.X(a[3]),.Y(b[3]),.Ci(c[2]));
full_adder a5(.Co(c[4]),.S(s[4]),.X(a[4]),.Y(b[4]),.Ci(c[3]));
full_adder a6(.Co(c[5]),.S(s[5]),.X(a[5]),.Y(b[5]),.Ci(c[4]));
full_adder a7(.Co(c[6]),.S(s[6]),.X(a[6]),.Y(b[6]),.Ci(c[5]));
full_adder a8(.Co(c[7]),.S(s[7]),.X(a[7]),.Y(b[7]),.Ci(c[6]));
full_adder a9(.Co(c[8]),.S(s[8]),.X(a[8]),.Y(b[8]),.Ci(c[7]));
full_adder a10(.Co(c[9]),.S(s[9]),.X(a[9]),.Y(b[9]),.Ci(c[8]));
full_adder a11(.Co(c[10]),.S(s[10]),.X(a[10]),.Y(b[10]),.Ci(c[9]));
full_adder a12(.Co(c[11]),.S(s[11]),.X(a[11]),.Y(b[11]),.Ci(c[10]));
full_adder a13(.Co(c[12]),.S(s[12]),.X(a[12]),.Y(b[12]),.Ci(c[11]));
full_adder a14(.Co(c[13]),.S(s[13]),.X(a[13]),.Y(b[13]),.Ci(c[12]));
full_adder a15(.Co(c[14]),.S(s[14]),.X(a[14]),.Y(b[14]),.Ci(c[13]));
full_adder a16(.Co(c[15]),.S(s[15]),.X(a[15]),.Y(b[15]),.Ci(c[14]));
full_adder a17(.Co(c[16]),.S(s[16]),.X(a[16]),.Y(b[16]),.Ci(c[15]));
full_adder a18(.Co(c[17]),.S(s[17]),.X(a[17]),.Y(b[17]),.Ci(c[16]));
full_adder a19(.Co(c[18]),.S(s[18]),.X(a[18]),.Y(b[18]),.Ci(c[17]));
full_adder a20(.Co(c[19]),.S(s[19]),.X(a[19]),.Y(b[19]),.Ci(c[18]));
full_adder a21(.Co(c[20]),.S(s[20]),.X(a[20]),.Y(b[20]),.Ci(c[19]));
full_adder a22(.Co(c[21]),.S(s[21]),.X(a[21]),.Y(b[21]),.Ci(c[20]));
full_adder a23(.Co(c[22]),.S(s[22]),.X(a[22]),.Y(b[22]),.Ci(c[21]));
full_adder a24(.Co(c[23]),.S(s[23]),.X(a[23]),.Y(b[23]),.Ci(c[22]));
full_adder a25(.Co(c[24]),.S(s[24]),.X(a[24]),.Y(b[24]),.Ci(c[23]));
full_adder a26(.Co(c[25]),.S(s[25]),.X(a[25]),.Y(b[25]),.Ci(c[24]));
full_adder a27(.Co(c[26]),.S(s[26]),.X(a[26]),.Y(b[26]),.Ci(c[25]));
full_adder a28(.Co(c[27]),.S(s[27]),.X(a[27]),.Y(b[27]),.Ci(c[26]));
full_adder a29(.Co(c[28]),.S(s[28]),.X(a[28]),.Y(b[28]),.Ci(c[27]));
full_adder a30(.Co(c[29]),.S(s[29]),.X(a[29]),.Y(b[29]),.Ci(c[28]));
full_adder a31(.Co(c[30]),.S(s[30]),.X(a[30]),.Y(b[30]),.Ci(c[29]));
full_adder a32(.Co(overflow),.S(s[31]),.X(a[31]),.Y(b[31]),.Ci(c[30]));
endmodule
